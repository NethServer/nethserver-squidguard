Unknown=
Title=F&ouml;rbjuden
Prefix=Access till denna sida &auml;r stoppad:
Suffix=
Info=Mer information om ufdbGuard &auml;r
Here=h&auml;r
